module example
fn main() {
	print("Hello World")
}
