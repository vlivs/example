module vlivs/example
func main() {
	print("Hello World")
}
