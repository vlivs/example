module example
func main() {
	print("Hello World")
}
